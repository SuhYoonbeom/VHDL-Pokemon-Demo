library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package torterra_pkg is
    ----------------------------------------------------------------
    -- Torterra sprite dimensions and types
    ----------------------------------------------------------------
    constant TORTERRA_W : integer := 80;
    constant TORTERRA_H : integer := 80;

    subtype tort_color_t is std_logic_vector(3 downto 0);
    type    tort_row_t    is array(0 to TORTERRA_W-1) of tort_color_t;
    type    tort_sprite_t is array(0 to TORTERRA_H-1) of tort_row_t;

    -- 80x80 color-index sprite (front-facing Torterra)
    constant TORTERRA_FRONT : tort_sprite_t;

    -- Color mapping for Torterra sprite
    procedure torterra_color(
        color_idx : in  std_logic_vector(3 downto 0);
        r_out     : out std_logic_vector(3 downto 0);
        g_out     : out std_logic_vector(3 downto 0);
        b_out     : out std_logic_vector(3 downto 0)
    );
end package torterra_pkg;

package body torterra_pkg is

    -- *** your big 80x80 array, just renamed ***
    constant TORTERRA_FRONT : tort_sprite_t := (
        -- row 0 ..
        0 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        1 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1101", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        2 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1101", "1100", "1100", "1100", "1101", "1101", "0000", "1101", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        3 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1101", "0000", "0000", "0000", "0000", "1101", "1101", "1100", "1100", "1011", "1011", "1100", "1100", "1100", "1101", "1100", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        4 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1100", "1011", "1100", "1101", "1101", "0000", "0000", "1101", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        5 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1011", "1100", "1011", "1011", "1011", "1100", "1101", "1101", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        6 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1101", "1100", "1100", "1011", "1011", "1011", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        7 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        8 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "1100", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        9 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "0000", "1101", "1101", "1101", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        10 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1100", "1100", "1011", "1011", "1011", "1011", "1100", "1011", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "1101", "1100", "1011", "1011", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        11 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1100", "1100", "1011", "1011", "1100", "1011", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "1101", "1101", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        12 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1101", "1011", "1011", "1011", "1011", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1101", "0000", "0000", "0000", "0000", "0000", "0000"),
        13 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1011", "1011", "1101", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1101", "1100", "1100", "0001", "0000", "0000", "0000", "0000", "0000", "0000"),
        14 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1011", "1011", "1101", "1101", "1011", "1011", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "0001", "0000", "0000", "0000", "0000", "0000", "0000"),
        15 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0011", "0000", "0000", "0000", "0000", "1101", "1100", "1011", "1011", "1011", "1100", "1100", "1100", "1011", "1011", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "1101", "1011", "1011", "1011", "1101", "1101", "1100", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        16 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0100", "0011", "0000", "0000", "0000", "0000", "1101", "1100", "1100", "1100", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1011", "1011", "1011", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        17 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0100", "0100", "0011", "0000", "0000", "0000", "0000", "0001", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "1000", "0001", "1101", "1101", "1101", "0001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "0001", "0000", "0000", "0000", "0000", "0000", "0000"),
        18 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0100", "0100", "0100", "0011", "0000", "0000", "0000", "0000", "0000", "0001", "1101", "1101", "1101", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1000", "0001", "1000", "1000", "0001", "1101", "1101", "1101", "0001", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1101", "0000", "0000", "0000", "0000", "0000", "0000"),
        19 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0101", "0100", "0100", "0100", "0100", "0011", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "1101", "1101", "1101", "1101", "1101", "0001", "1101", "0001", "0001", "1000", "1000", "1000", "1000", "1101", "1101", "0001", "0001", "1100", "1100", "1100", "1011", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1011", "1100", "1011", "1011", "1011", "1011", "1101", "0000", "0000", "0000", "0000", "0000"),
        20 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0001", "0000", "0000", "0000", "0011", "0100", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0001", "1000", "1000", "0001", "1101", "1101", "0001", "1100", "1100", "1100", "1101", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1100", "1011", "1100", "1011", "1011", "1100", "1100", "0001", "0000", "0000", "0000", "0000"),
        21 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0100", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0001", "0000", "0000", "0100", "0100", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "1000", "1000", "1000", "1101", "1101", "0001", "1100", "1100", "0001", "1101", "0001", "0001", "1100", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1100", "1100", "0001", "0000", "0000", "0000", "0000"),
        22 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0001", "0000", "0011", "0100", "0100", "0100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "1000", "0110", "0110", "0001", "1101", "1101", "0001", "0001", "1100", "0001", "1000", "0110", "0001", "0001", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "0001", "0000", "0000", "0000", "0000"),
        23 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0011", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "1100", "1100", "0001", "0011", "0100", "0100", "0100", "1101", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1000", "0110", "0110", "0001", "1101", "1101", "1101", "1101", "1000", "1000", "0110", "0110", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "0001", "0000", "0000", "0000", "0000", "0000"),
        24 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0100", "0011", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "1100", "1100", "1100", "1100", "1100", "0001", "0100", "0100", "0100", "0100", "0011", "0001", "0001", "1101", "1101", "0001", "0001", "1101", "1101", "1101", "0001", "1101", "1000", "0110", "0110", "0110", "0001", "1101", "1000", "1000", "0110", "0110", "0110", "1000", "1000", "0001", "0001", "1100", "1100", "0001", "0001", "0001", "1101", "1100", "1100", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000"),
        25 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0100", "0100", "0011", "0000", "0000", "0000", "0011", "0100", "0101", "0101", "0101", "0011", "1100", "1011", "1100", "1100", "1100", "1100", "0001", "0100", "0100", "0100", "0100", "0011", "0011", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0000", "0001", "0110", "0111", "0111", "0110", "1000", "0110", "0111", "0111", "0110", "1000", "1000", "1101", "1101", "1101", "1101", "0001", "0001", "1101", "0001", "0000", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        26 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0100", "0100", "0011", "0000", "0000", "1100", "1100", "1100", "0100", "0100", "0011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "0001", "0100", "0100", "0100", "0011", "0011", "0011", "0011", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0111", "0111", "1000", "0111", "0111", "0111", "0110", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        27 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0100", "0100", "0100", "0011", "1001", "1100", "1011", "1011", "1100", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0011", "0011", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "1000", "0111", "0111", "0110", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        28 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0100", "0100", "0100", "0100", "1001", "1011", "1011", "1011", "1011", "1011", "1100", "1001", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0001", "1000", "1000", "1000", "1000", "1000", "0000", "1000", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "1000", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        29 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "1001", "1011", "1100", "1100", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "0110", "0110", "0110", "1000", "1000", "0111", "0111", "1000", "0110", "0110", "1000", "1000", "0110", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        30 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "1001", "1011", "1011", "1100", "1100", "1100", "1001", "1001", "1001", "1001", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1000", "1000", "0111", "0111", "1000", "1000", "1000", "1000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0001", "0001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        31 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "1100", "1100", "1100", "1100", "1100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1000", "0111", "0111", "1000", "1000", "0110", "0110", "0110", "1000", "0110", "0110", "1000", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0001", "0001", "1101", "1101", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        32 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "1001", "1011", "1011", "1100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1011", "1011", "1000", "1000", "0110", "0111", "1000", "0110", "0110", "0001", "0001", "0001", "1000", "0110", "0110", "1000", "0110", "0110", "1000", "0001", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        33 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0100", "0100", "1001", "1001", "1011", "1100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1000", "0111", "0111", "0111", "0111", "0001", "0001", "1001", "1001", "1100", "1100", "1001", "1001", "1000", "0110", "0110", "0110", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        34 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1001", "1001", "1011", "1011", "1100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "1001", "1000", "0111", "1000", "0001", "0001", "1001", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1000", "0110", "0111", "0111", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        35 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1011", "1011", "1011", "1011", "1011", "1100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "1001", "1000", "1000", "1001", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1001", "1000", "0111", "0111", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        36 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1001", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1000", "0111", "0110", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        37 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1001", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1000", "0111", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        38 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1011", "1011", "1011", "1011", "1011", "1001", "1001", "1001", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0110", "0111", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0001", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        39 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "1011", "1011", "1011", "1001", "1001", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "0111", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        40 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1001", "1001", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "0110", "1000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        41 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0111", "0111", "1011", "1011", "0111", "0111", "0111", "0111", "0111", "1000", "0110", "1000", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1001", "1010", "1010", "1001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        42 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0111", "0111", "0111", "0111", "0110", "1000", "0110", "0110", "0001", "0001", "0000", "0000", "0000", "0000", "1001", "1010", "1010", "1010", "1010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        43 => ("0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0101", "0001", "0000", "0000", "1001", "1001", "1001", "1001", "1010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        44 => ("0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0001", "0001", "0001", "0001", "1010", "1010", "1010", "1010", "1010", "1010", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0101", "0100", "0001", "1001", "1010", "1010", "1010", "1010", "1001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        45 => ("0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0100", "0100", "0100", "0011", "0001", "0001", "1010", "1010", "1001", "1010", "1010", "1011", "1011", "1011", "1011", "1010", "1010", "1010", "1010", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0001", "0101", "0100", "0001", "1010", "1010", "1010", "1010", "1010", "1001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        46 => ("0000", "0000", "0000", "0000", "0000", "0000", "0011", "0101", "0100", "0011", "0001", "0001", "1010", "1010", "1010", "1001", "1010", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "1010", "1010", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1001", "1001", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "1001", "1001", "1001", "0110", "0101", "0101", "0100", "0001", "1001", "1001", "1010", "1010", "1010", "1010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        47 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0011", "0011", "0010", "0001", "1010", "1010", "1010", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "1010", "0001", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0001", "1010", "1010", "1001", "1010", "1010", "1010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        48 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "1010", "1010", "1001", "1011", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "1010", "0001", "1010", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0001", "1010", "1010", "1010", "1010", "1001", "1010", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        49 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0010", "1001", "1011", "1001", "1010", "1011", "1011", "1011", "1011", "1011", "1010", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "1010", "0001", "1010", "1010", "1010", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0001", "0001", "1010", "1010", "1010", "1010", "1001", "1010", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        50 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0010", "0010", "0101", "0101", "1001", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "0010", "0010", "0010", "1010", "1010", "1010", "1010", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0001", "0001", "0001", "1010", "0001", "1010", "1010", "1010", "1010", "1010", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        51 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0010", "0010", "1011", "1011", "1011", "1010", "1001", "1010", "0101", "0101", "0010", "0010", "0010", "1010", "1010", "1010", "1010", "0001", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0001", "0001", "0001", "1010", "1010", "1010", "1010", "0001", "1010", "1010", "1010", "0110", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        52 => ("0000", "0000", "0000", "0000", "0000", "0000", "0001", "0100", "0100", "0101", "0101", "0101", "0101", "1001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0010", "0101", "0010", "1011", "1011", "1011", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0010", "0010", "1010", "1010", "1010", "1010", "1010", "1010", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "1010", "1010", "1010", "1001", "1000", "1000", "0001", "1010", "1010", "0110", "0110", "0110", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        53 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0100", "0100", "0100", "0100", "0001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "0010", "0110", "0101", "0001", "1011", "1010", "1001", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0010", "0010", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1010", "1010", "1010", "1000", "1000", "0110", "0110", "1000", "0110", "0110", "0110", "0111", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        54 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0100", "0100", "0001", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "0010", "0101", "0101", "0100", "0001", "1010", "1010", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1010", "1010", "1000", "1000", "0110", "0110", "0110", "0110", "0001", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        55 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0001", "0001", "0001", "1011", "0010", "0010", "0010", "0010", "0010", "0010", "1010", "0010", "0001", "0010", "0100", "0010", "0010", "1000", "1001", "1001", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0001", "0001", "1011", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1010", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        56 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0110", "0110", "0001", "0010", "0011", "0011", "0011", "0011", "0011", "0011", "0010", "0111", "0111", "0001", "0001", "0001", "0111", "1000", "1010", "1010", "1001", "1001", "0100", "0100", "0100", "0001", "0001", "0001", "0001", "1011", "1011", "1011", "1011", "1011", "1011", "1000", "1000", "1000", "1000", "1010", "1010", "1010", "1010", "1010", "1001", "1010", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        57 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0110", "0110", "0110", "0001", "0010", "0011", "0011", "0011", "0011", "0011", "0010", "0001", "0111", "0111", "0111", "0111", "0111", "1000", "1000", "1010", "1010", "1010", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "1010", "1011", "1011", "1011", "1011", "1000", "1000", "0111", "0111", "0111", "0111", "1000", "1010", "1010", "1010", "1010", "1001", "1010", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        58 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0010", "0011", "0011", "0011", "0010", "0010", "0001", "0111", "0111", "1000", "1001", "1000", "1010", "1010", "1010", "1010", "1001", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "1010", "0001", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "1000", "1010", "1010", "1000", "1001", "1000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        59 => ("0000", "0000", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0010", "0010", "0010", "0010", "0001", "0010", "0001", "1000", "1000", "1000", "1010", "1010", "1010", "1010", "1001", "1001", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0001", "1000", "1000", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        60 => ("0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "1000", "0001", "0010", "0010", "0010", "0010", "0010", "0001", "1010", "1010", "1010", "1010", "1001", "0001", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "1000", "0110", "0110", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        61 => ("0000", "0000", "0000", "0000", "0000", "1000", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0010", "0010", "0010", "0001", "1001", "1001", "1001", "0001", "0001", "0001", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0001", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        62 => ("0000", "0000", "0000", "0000", "0000", "1000", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0010", "0010", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0001", "0110", "0110", "0110", "0001", "0110", "0110", "0110", "0110", "0110", "1000", "0110", "0110", "0110", "0110", "0110", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        63 => ("0000", "0000", "0000", "0000", "0000", "1000", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "1000", "1000", "1000", "0110", "0110", "1000", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "1000", "1000", "0001", "0001", "0000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        64 => ("0000", "0000", "0000", "0000", "0000", "1000", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "1000", "1000", "1000", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0001", "0000", "0000", "0000", "0001", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        65 => ("0000", "0000", "0000", "0000", "1000", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0110", "0110", "0110", "0110", "0110", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "1000", "0110", "0110", "0110", "0110", "0110", "1000", "0100", "0011", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        66 => ("0000", "0000", "0000", "0000", "1000", "0111", "1000", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "1000", "0111", "0111", "0111", "0111", "1000", "0111", "0111", "0111", "0111", "0111", "1000", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0001", "0110", "1000", "0110", "0110", "1000", "0100", "0100", "0100", "1000", "1000", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        67 => ("0000", "0000", "0000", "0000", "0010", "0011", "0101", "0101", "0010", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0001", "1000", "0100", "0110", "0110", "1000", "0100", "0100", "0100", "1000", "0100", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        68 => ("0000", "0000", "0000", "0000", "0010", "0011", "0101", "0101", "0100", "0010", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0111", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0001", "1000", "0100", "1000", "1000", "0100", "0100", "0100", "0100", "0010", "0100", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        69 => ("0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0010", "0110", "0110", "1000", "0100", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0010", "0100", "0100", "1000", "0100", "0100", "0100", "0100", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        70 => ("0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0110", "1000", "0100", "0100", "0100", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        71 => ("0000", "0000", "0000", "0000", "0011", "0101", "0101", "0101", "0100", "0100", "0110", "1000", "0100", "0100", "0100", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0011", "0101", "0011", "0110", "0110", "0110", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        72 => ("0000", "0000", "0000", "0000", "0011", "0101", "0101", "0100", "0100", "0010", "0001", "0001", "0010", "0010", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0110", "0111", "0111", "0111", "0110", "0011", "0101", "0101", "0101", "0011", "0110", "0100", "1000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        73 => ("0000", "0000", "0000", "0000", "0000", "0010", "0010", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0011", "0011", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0100", "0110", "0100", "0100", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        74 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0101", "0101", "0110", "0110", "0011", "0101", "0101", "0101", "0101", "0100", "0110", "0100", "0100", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        75 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0101", "0101", "0011", "0110", "0011", "0101", "0101", "0101", "0101", "0100", "0010", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        76 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0010", "0001", "0001", "0001", "0001", "0100", "0100", "0100", "0100", "0100", "0010", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        77 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0010", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        78 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000"),
        79 => ("0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000")
    );

    ----------------------------------------------------------------
    -- Torterra color mapping (using provided palette)
    ----------------------------------------------------------------
    procedure torterra_color(
        color_idx : in  std_logic_vector(3 downto 0);
        r_out     : out std_logic_vector(3 downto 0);
        g_out     : out std_logic_vector(3 downto 0);
        b_out     : out std_logic_vector(3 downto 0)
    ) is
    begin
        case color_idx is
            when "0000" =>  -- 0: transparent / black
                r_out := "0000";
                g_out := "0000";
                b_out := "0000";

            when "0001" =>  -- 1: #282828
                r_out := "0010";
                g_out := "0010";
                b_out := "0010";

            when "0010" =>  -- 2: #485058
                r_out := "0100";
                g_out := "0101";
                b_out := "0101";

            when "0011" =>  -- 3: #687078
                r_out := "0110";
                g_out := "0111";
                b_out := "0111";

            when "0100" =>  -- 4: #B8B8B8
                r_out := "1011";
                g_out := "1011";
                b_out := "1011";

            when "0101" =>  -- 5: #E0E0E0
                r_out := "1110";
                g_out := "1110";
                b_out := "1110";

            when "0110" =>  -- 6: #886840
                r_out := "1000";
                g_out := "0110";
                b_out := "0100";

            when "0111" =>  -- 7: #B08051
                r_out := "1011";
                g_out := "1000";
                b_out := "0101";

            when "1000" =>  -- 8: #614837
                r_out := "0110";
                g_out := "0100";
                b_out := "0011";

            when "1001" =>  -- 9: #385828
                r_out := "0011";
                g_out := "0101";  -- if you had "0101" here before, keep it
                b_out := "0010";

            when "1010" =>  -- 10: #587841
                r_out := "0101";
                g_out := "0111";
                b_out := "0100";

            when "1011" =>  -- 11: #40A840
                r_out := "0100";
                g_out := "1010";
                b_out := "0100";

            when "1100" =>  -- 12: #308838
                r_out := "0011";
                g_out := "1000";
                b_out := "0011";

            when "1101" =>  -- 13: #186018
                r_out := "0001";
                g_out := "0110";
                b_out := "0001";

            -- 14, 15 are unused -> treat as transparent/black
            when others =>
                r_out := "0000";
                g_out := "0000";
                b_out := "0000";
        end case;
    end procedure torterra_color;

end package body torterra_pkg;
