library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity alphabet is
    port (
        char_code : in  std_logic_vector(5 downto 0); -- 0-9, A-Z
        glyph_x   : in  std_logic_vector(2 downto 0); -- 0..4
        glyph_y   : in  std_logic_vector(2 downto 0); -- 0..6
        pixel_on  : out std_logic                     -- '1' = draw
    );
end entity alphabet;

architecture Behavioral of alphabet is

    subtype row_t   is std_logic_vector(4 downto 0);  -- 5 columns
    type    glyph_t is array(0 to 6) of row_t;        -- 7 rows
    type    font_t  is array(0 to 35) of glyph_t;     -- 0-9, A-Z

    -- 5x7 font:
    -- index 0-9   : '0'..'9'
    -- index 10-35 : 'A'..'Z'
    constant FONT : font_t := (
         0 => ("01110","10001","10011","10101","11001","10001","01110"), -- '0'
         1 => ("00100","01100","00100","00100","00100","00100","01110"), -- '1'
         2 => ("01110","10001","00001","00010","00100","01000","11111"), -- '2'
         3 => ("01110","10001","00001","00110","00001","10001","01110"), -- '3'
         4 => ("00010","00110","01010","10010","11111","00010","00010"), -- '4'
         5 => ("11111","10000","11110","00001","00001","10001","01110"), -- '5'
         6 => ("01110","10000","11110","10001","10001","10001","01110"), -- '6'
         7 => ("11111","00001","00010","00100","01000","01000","01000"), -- '7'
         8 => ("01110","10001","10001","01110","10001","10001","01110"), -- '8'
         9 => ("01110","10001","10001","01111","00001","00010","01100"), -- '9'
        10 => ("01110","10001","10001","11111","10001","10001","10001"), -- 'A'
        11 => ("11110","10001","10001","11110","10001","10001","11110"), -- 'B'
        12 => ("01110","10001","10000","10000","10000","10001","01110"), -- 'C'
        13 => ("11100","10010","10001","10001","10001","10010","11100"), -- 'D'
        14 => ("11111","10000","10000","11110","10000","10000","11111"), -- 'E'
        15 => ("11111","10000","10000","11110","10000","10000","10000"), -- 'F'
        16 => ("01110","10001","10000","10000","10011","10001","01110"), -- 'G'
        17 => ("10001","10001","10001","11111","10001","10001","10001"), -- 'H'
        18 => ("11111","00100","00100","00100","00100","00100","11111"), -- 'I'
        19 => ("00001","00001","00001","00001","10001","10001","01110"), -- 'J'
        20 => ("10001","10010","10100","11000","10100","10010","10001"), -- 'K'
        21 => ("10000","10000","10000","10000","10000","10000","11111"), -- 'L'
        22 => ("10001","11011","10101","10101","10001","10001","10001"), -- 'M'
        23 => ("10001","11001","10101","10011","10001","10001","10001"), -- 'N'
        24 => ("01110","10001","10001","10001","10001","10001","01110"), -- 'O'
        25 => ("11110","10001","10001","11110","10000","10000","10000"), -- 'P'
        26 => ("01110","10001","10001","10001","10101","10010","01101"), -- 'Q'
        27 => ("11110","10001","10001","11110","10100","10010","10001"), -- 'R'
        28 => ("01111","10000","10000","01110","00001","00001","11110"), -- 'S'
        29 => ("11111","00100","00100","00100","00100","00100","00100"), -- 'T'
        30 => ("10001","10001","10001","10001","10001","10001","01110"), -- 'U'
        31 => ("10001","10001","10001","10001","10001","01010","00100"), -- 'V'
        32 => ("10001","10001","10001","10101","10101","11011","10001"), -- 'W'
        33 => ("10001","10001","01010","00100","01010","10001","10001"), -- 'X'
        34 => ("10001","10001","01010","00100","00100","00100","00100"), -- 'Y'
        35 => ("11111","00001","00010","00100","01000","10000","11111")  -- 'Z'
    );

begin
    process(char_code, glyph_x, glyph_y)
        variable x, y   : integer;
        variable idx    : integer;
        variable on_v   : std_logic;
        variable bitpos : integer;
    begin
        x   := to_integer(unsigned(glyph_x)); -- 0..4
        y   := to_integer(unsigned(glyph_y)); -- 0..6
        idx := to_integer(unsigned(char_code));
        on_v := '0';

        if (idx >= 0 and idx <= 35) and
           (x >= 0 and x <= 4) and
           (y >= 0 and y <= 6) then
            -- row y, column x (leftmost bit is index 4)
            bitpos := 4 - x;
            if FONT(idx)(y)(bitpos) = '1' then
                on_v := '1';
            end if;
        else
            on_v := '0';
        end if;

        pixel_on <= on_v;
    end process;

end architecture Behavioral;
